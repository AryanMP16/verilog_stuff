//module register_file (input [5 : 0] read_address/*if msb = 1, read data; otherwise RT*/, input [4 : 0] write_address, input [15 : 0] data_in);
	